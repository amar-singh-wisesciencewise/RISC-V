


`timescale 1ns / 1ps


// This module combine RISC V CPU and Instruction and Data memory

module risc_v_microcontroller();

//instantiate RISC V CPU; IMEM and DMEM.




endmodule
